

module adder(adder_if.dut_md inf);
  
  // addition operation
  assign inf.s = inf.a + inf.b;

endmodule
